module gate_level(a,b,c);
  input a,b;
  output c;
  and(c,a,b);
endmodule
